typedef enum {TRANS, RECEIVE, REPEATER} tr_type;

class Transaction;
    bit [31:0] data;
    int id;
endclass

module class_example;
    Transaction tr[tr_type]; // asociativo
    
    initial begin
        tr[TRANS]    = new();
        tr[RECEIVE]  = new();
        tr[REPEATER] = new();

        foreach(tr[i]) begin 
          tr[i].data = i*i;
          tr[i].id = i+1;
        end

        foreach(tr[i]) $display("tr[%0s].data = %0d, tr[%0s].id = %0d",i.name, tr[i].data, i.name, tr[i].id);
    end
endmodule